/* Copyright 2023 Fereie

   Licensed under the Apache License, Version 2.0 (the "License");
   you may not use this file except in compliance with the License.
   You may obtain a copy of the License at

       http://www.apache.org/licenses/LICENSE-2.0

   Unless required by applicable law or agreed to in writing, software
   distributed under the License is distributed on an "AS IS" BASIS,
   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
   See the License for the specific language governing permissions and
   limitations under the License.
*/

// 2 flip flop synchonizer
`timescale 1ns / 1ps

module doubleff_sync(clk,rst,d,q);
parameter WIDTH = 4;

input clk,rst;
input [WIDTH-1:0] d;
output reg [WIDTH-1:0] q;
reg [WIDTH-1:0] d1d2_0;

always @(posedge clk or negedge rst) begin
   if(!rst) begin
     {d1d2_0,q} <= 0;
   end
   else begin
       d1d2_0 <= d;
       q <= d1d2_0;
       end
end


endmodule
